-- This is the top level file for the SAP-1 project

library ieee;
use ieee.std_logic_1164.all;

entity sap_1_top is
    port (
        i_Ext_Clk : in std_logic
    );
end entity sap_1_top;

architecture  rtl of sap_1_top is
begin
end rtl;